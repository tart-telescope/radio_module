module ser_pll(input clkin, output clkout);

endmodule
